library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

entity ALU is
  port(
    src1, src2: in STD_LOGIC_VECTOR(31 downto 0);
    ALUcontrol: in STD_LOGIC_VECTOR(2 downto 0);
    result: out STD_LOGIC_VECTOR(31 downto 0);
    zero: out std_logic
  );
end ALU;

architecture behav of ALU is
signal res_buff : STD_LOGIC_VECTOR(31 downto 0);
begin
  process(ALUcontrol) 
    begin
    case ALUcontrol is
      when "000" => res_buff <= (src1 AND src2);
      when "001" => res_buff <= (src1 or src2);
      when "010" => res_buff <= (src1 + src2);
      when "100" => res_buff <= (src1 AND NOT src2);
      when "101" => res_buff <= (src1 OR NOT src2);
      when "110" => res_buff <= (src1 - src2);
      when "111" =>
        if(src1 < src2) then
          res_buff <= "00000000000000000000000000000001";
        else
          res_buff <= "00000000000000000000000000000000";
        end if;
      when others => NULL;
    end case;

    if res_buff = 0 then
      zero <= '1';
    else
      zero <= '0';
    end if;
  result <= res_buff;
  end process;
end behav;
 
