library ieee;
use ieee.std_logic_1164.all;

entity shiftleft2_32b is
  Port(
    A: in STD_LOGIC_VECTOR(31 downto 0);
    Z: out STD_LOGIC_VECTOR(31 downto 0)
  );
end;

architecture behav of shiftleft2_32b is
  begin
    Z <= A(29 downto 0) & "00";
end;
