library ieee;
use ieee.std_logic_1164.all;

entity shiftleft2_26b is
  Port(
    A: in STD_LOGIC_VECTOR(25 downto 0);
    Z: out STD_LOGIC_VECTOR(27 downto 0)
  );
end ;
architecture behav of shiftleft2_26b is
  begin
    Z <= A & "00";
end;
